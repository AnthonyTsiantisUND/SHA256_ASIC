module SHA256 #() (
	input logic clk, reset,
	input logic[15:0] input_data,
	output logic[15:0] encrypted_data
);



endmodule
